class ddr3_tb_driver extends uvm_driver;
    function new();
        
    endfunction //new()
endclass //ddr3_tb_driver extends uvm_drive