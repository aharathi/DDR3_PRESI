/// testbench components ///
